library ieee;
use ieee.std_logic_1164.all;


package State_Package is

	-- Definition of variable for a finite state machine
   TYPE State_type IS (GREENS, YELLOWS, REDS);  -- Define the states
   
end package State_Package;