library ieee;
use ieee.std_logic_1164.all;
 
package State_Package is
 
   TYPE State_type IS (GREENS, YELLOWS, REDS);  -- Define the states
   
end package State_Package;